module LOSUJ(KEY, HEX0);


endmodule