//Zadanie 1
module LOSOWE